//============================================================================//
//                                                                            //
//      Parameterize Wishbone Slave Template                                  //
//                                                                            //
//      Module name: wbs_template                                             //
//      Desc: parameterized wishbone slave template, with byte enables and    //
//            parameterized address and data widths.                          //
//      Date: July 2012                                                       //
//      Developer: Wesley New                                                 //
//      Licence: GNU General Public License ver 3                             //
//      Notes:                                                                //
//                                                                            //
//============================================================================//

module wbs_template #(
      //=============
      // parameters
      //=============
      parameter DEV_BASE_ADDR  = {BUS_ADDR_WIDTH{1'b0}}, // default 32'h0
      parameter DEV_HIGH_ADDR  = {{(BUS_ADDR_WIDTH-4){1'b0}}, 4'hF}, // default 32'h000000EE
      parameter BUS_DATA_WIDTH = 32,  // default is 32. but can be 8, 16, 32, 64
      parameter BUS_ADDR_WIDTH = 8    // default is 8.  but can be 4, 8, 16, 32
   ) (
      //===============
      // fabric ports
      //===============
      input        fabric_clk,
      input [31:0] fabric_data_in,
      
      //============
      // wb inputs
      //============
      input                      wb_clk_i,
      input                      wb_rst_i,
      input                      wbs_cyc_i,
      input                      wbs_stb_i,
      input                      wbs_we_i,
      input  [BYTE_EN_WIDTH-1:0] wbs_sel_i,
      input [BUS_ADDR_WIDTH-1:0] wbs_adr_i,
      input [BUS_DATA_WIDTH-1:0] wbs_dat_i,
      
      //=============
      // wb outputs
      //=============
      output reg [BUS_DATA_WIDTH-1:0] wbs_dat_o,
      output reg                      wbs_ack_o,
      output reg                      wbs_err_o,
      output reg                      wbs_int_o
   );
   
   //===================
   // local parameters
   //===================
   // byte enable is always the data width/8
   // thus the data width is only able to be multiples of 8
   localparam BYTE_EN_WIDTH = BUS_DATA_WIDTH / 8;
   
   //========
   // wires
   //========
   wire adr_match = wbs_adr_i >= DEV_BASE_ADDR && wbs_adr_i <= DEV_HIGH_ADDR;

   //============
   // registers
   //============
   reg [BUS_DATA_WIDTH-1:0] reg_buf_i = {BUS_DATA_WIDTH{1'b0}};

   //blocks
   always @ (posedge wb_clk_i) begin
      // reset logic
      if (wb_rst_i) begin
         wbs_dat_o <= {BUS_DATA_WIDTH{1'b0}};
         wbs_ack_o <= 0;
         wbs_int_o <= 0;
      end
   
      else begin
         // when the master acks our ack, then put our ack down
         if (wbs_ack_o & ~wbs_stb_i) begin
            wbs_ack_o <= 0;
         end
         // master is requesting somethign
         if (adr_match & wbs_stb_i & wbs_cyc_i) begin
            //================
            // write request
            //================
            if (wbs_we_i) begin
               // bring the address down to the base address
               case (wbs_adr_i - DEV_BASE_ADDR)
                  // writing something to address
                  32'h0: begin
                     // byte enabled writes
                     if (wbs_sel_i[0])
                        reg_buf_i  [7:0] <= wbs_dat_i[7:0];
                     if (wbs_sel_i[1])
                        reg_buf_i [15:8] <= wbs_dat_i[15:8];
                     if (wbs_sel_i[2])
                        reg_buf_i[23:16] <= wbs_dat_i[23:16];
                     if (wbs_sel_i[3])
                        reg_buf_i[31:24] <= wbs_dat_i[31:24];
   
                     $display("user wrote %h", reg_buf_i);
                  end
                  //add as many addresses as you need here
                  default: begin
                     $display("no case for write address %h", wbs_adr_i);
                  end
               endcase
            end
            
            //===============
            // read request
            //===============
            else begin 
               case (wbs_adr_i)
                  32'h0: begin
                     //reading something from address 0
                     $display("user read %h", reg_buf_i);
                     wbs_dat_o <= reg_buf_i;
                  end
                  //add as many addresses as you need here
                  default: begin
                     $display("no case for read address %h", wbs_adr_i);
                  end
               endcase
            end
            wbs_ack_o <= 1;
         end
      end
   end
endmodule
